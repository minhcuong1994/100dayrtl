interface alu_interface (input clk);
  logic rst_n;
  logic [2:0] ctl;
  logic [7:0]a, b, q;
  logic cout;
  
  
endinterface