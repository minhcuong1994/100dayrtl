`timescale 1ns/1ns

`define PARITY_EVEN

//compare output dut vs. model task ---------------------------------------------
task compare;
  input [7:0]dut_out;
  input dut_done;
  input dut_err;
  
  input [7:0] mdl_out;
  input mdl_done;
  input mdl_err;
    
  if ((mdl_done != dut_done) | (mdl_out != dut_out) | (mdl_err != dut_err)) begin
    $display("ERROR! mdl_done=%b, mdl_out=%b, mdl_err=%b, dut_done=%b, dut_out=%b, dut_err=%b",mdl_done, mdl_out, mdl_err, dut_done, dut_out, dut_err);
  end else
    $display("PASS");

endtask


//parity calculator func---------------------------------------------------------
function logic parity_cal(input [7:0] data);
  
  logic [4:0] p_sum;
  
  p_sum = data[0] + data[1] + data[2] + data[3] + data[4] + data[5] + data[6];
  
  `ifdef PARITY_EVEN
  if ((p_sum % 2) != data[7]) parity_cal = 1'b1;
  else parity_cal = 1'b0;
  `endif
  
  `ifdef PARITY_ODD
  if (((p_sum + 1)% 2) != data[7]) parity_cal = 1'b1;
  else parity_cal = 1'b0;
  `endif
  
endfunction


//Testbench ---------------------------------------------------------------------
module testbench ();
  logic clk;
  logic rst_n, in;
  
  //signal get from dut
  logic [7:0] dut_out;
  logic dut_done;
  logic dut_err;
  
  //signal generated by model
  logic [7:0] mdl_out, mdl_out_temp;
  logic mdl_done;
  logic mdl_err;
  
  serial_rx dut(.clk(clk),
                .rst_n(rst_n),
                .in(in),
                .out(dut_out),
                .done(dut_done),
                .err(dut_err)
               );
  
  
  //clock initial
  initial begin 
    clk = 0;
  end
  always @ * begin
    clk <= #1 ~clk;
  end
  
  
  //simulation
  initial begin
    $dumpfile("file.vcd");
    $dumpvars();
    
    #220;
    $finish();
    
  end
  
  //stimulus signal to dut
  initial begin
    
    repeat(3) begin
    
      //clear model vars
      mdl_done = 0;
      mdl_out = 8'd0;
      mdl_err = 0;

      //reset
      in = 1;
      rst_n = 0;

      //clear reset (IDLE)
      @(posedge clk);
      rst_n = 1;

      //START
      @(posedge clk);
      in = 0;

      //Transmit 8 bits data
      for(int i = 0; i<8; i++) begin
        @(posedge clk);
        in = $urandom_range(0,1);
        mdl_out_temp = {in, mdl_out_temp[7:1]};
      end

      //STOP
      @(posedge clk);
      in = 1;

      //START AGAIN (DONE)
      @(posedge clk);
      in = 0;
      mdl_done = 1;
      mdl_out = {0, mdl_out_temp[6:0]};
      mdl_err = parity_cal(mdl_out_temp);

      //TRANSMIT NEXT 1 bit
      @(posedge clk);
      in = $urandom_range(0,1);
      mdl_out_temp = {in, mdl_out_temp[7:1]};
      mdl_done = 0;
      mdl_err = 0;

      //Transmit next 7 bits
      for(int i = 0; i<7; i++) begin
        @(posedge clk);
        in = $urandom_range(0,1);
        mdl_out_temp = {in, mdl_out_temp[7:1]};
      end

      //STOP
      @(posedge clk);
      in = 1;

      //DONE (IDLE)
      @(posedge clk);
      in = 1;
      mdl_done = 1; 
      mdl_out = {0, mdl_out_temp[6:0]};
      mdl_err = parity_cal(mdl_out_temp);

      //IDLE
      @(posedge clk);
      in = 1;
      mdl_done = 0;
      mdl_err = 0;

      //START
      @(posedge clk);
      in = 0;

      //Transmit 8 bits data
      for(int i = 0; i<8; i++) begin
        @(posedge clk);
        in = $urandom_range(0,1);
        mdl_out_temp = {in, mdl_out_temp[7:1]};
      end

      //STOP
      @(posedge clk);
      in = 1;


      //DONE (IDLE)
      @(posedge clk);
      in = 1;
      mdl_done = 1;
      mdl_out = {0, mdl_out_temp[6:0]};
      mdl_err = parity_cal(mdl_out_temp);

      //IDLE
      @(posedge clk);
      in = 1;
      mdl_done = 0;
      mdl_err = 0;
    end   
  end
  
  //compare result
  always @(posedge mdl_done) begin
    compare(dut_out, dut_done, dut_err, mdl_out, mdl_done, mdl_err);
  end
  
endmodule



